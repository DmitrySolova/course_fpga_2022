library verilog;
use verilog.vl_types.all;
entity course_3_mult_vlg_vec_tst is
end course_3_mult_vlg_vec_tst;
